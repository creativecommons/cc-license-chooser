function cc_js_t(s) {
		 if (s == "Brazil") { return "Brasilien"; } 
 if (s == "Canada") { return "Kanada"; } 
 if (s == "Italy") { return "Italien"; } 
 if (s == "Creative Commons") { return "Creative Commons"; } 
 if (s == "Serbia") { return "Serbien"; } 
 if (s == "Malta") { return "Malta"; } 
 if (s == "France") { return "Frankrike"; } 
 if (s == "Peru") { return "Peru"; } 
 if (s == "Argentina") { return "Argentina"; } 
 if (s == "Norway") { return "Norway"; } 
 if (s == "New Zealand") { return "Nya Zeeland"; } 
 if (s == "Ecuador") { return "Ecuador"; } 
 if (s == "Czech Republic") { return "Tjeckien"; } 
 if (s == "Israel") { return "Israel"; } 
 if (s == "Australia") { return "Australien"; } 
 if (s == "Korea") { return "Korea"; } 
 if (s == "Singapore") { return "Singapore"; } 
 if (s == "Thailand") { return "Thailand"; } 
 if (s == "South Africa") { return "Sydafrika"; } 
 if (s == "We have updated the version of your license to the most recent one available.") { return "We have updated the version of your license to the most recent one available."; } 
 if (s == "Slovenia") { return "Slovenien"; } 
 if (s == "Guatemala") { return "Guatemala"; } 
 if (s == "The licensor permits others to copy, distribute and transmit the work. In return, licensees may not use the work for commercial purposes — unless they get the licensor's permission.") { return "Licensgivaren tillåter andra att kopiera, distribuera och sända verket. I gengäld får licenstagarna inte använda verket för kommersiella ändamål -- om de inte får licensgivarens tillstånd."; } 
 if (s == "Noncommercial") { return "Ickekommersiell"; } 
 if (s == "Puerto Rico") { return "Puerto Rico"; } 
 if (s == "Belgium") { return "Belgien"; } 
 if (s == "Germany") { return "Tyskland"; } 
 if (s == "We have updated the version of your license to the most recent one available in your jurisdiction.") { return "We have updated the version of your license to the most recent one available in your jurisdiction."; } 
 if (s == "Hong Kong") { return "Hong Kong"; } 
 if (s == "Poland") { return "Polen"; } 
 if (s == "Spain") { return "Spanien"; } 
 if (s == "This ${work_type} is licensed under a <a rel=\"license\" href=\"${license_url}\">Creative Commons ${license_name} License</a>.") { return "Detta ${work_type} är licensierat under en <a rel=\"license\" href=\"${license_url}\">Creative Commons ${license_name} Licens</a>."; } 
 if (s == "Remix") { return "Remix"; } 
 if (s == "Netherlands") { return "Nederländerna"; } 
 if (s == "UK: England & Wales") { return "UK: England & Wales"; } 
 if (s == "Chile") { return "Chile"; } 
 if (s == "Unported") { return "Unported"; } 
 if (s == "Denmark") { return "Danmark"; } 
 if (s == "Philippines") { return "Filippinerna"; } 
 if (s == "Finland") { return "Finland"; } 
 if (s == "Macedonia") { return "Makedonien"; } 
 if (s == "United States") { return "Förenta Staterna"; } 
 if (s == "Sweden") { return "Sverige"; } 
 if (s == "No license chosen") { return "No license chosen"; } 
 if (s == "Croatia") { return "Kroatien"; } 
 if (s == "Luxembourg") { return "Luxemburg"; } 
 if (s == "Japan") { return "Japan"; } 
 if (s == "Switzerland") { return "Schweiz"; } 
 if (s == "UK: Scotland") { return "UK: Skottland"; } 
 if (s == "With a Creative Commons license, you keep your copyright but allow people to copy and distribute your work provided they give you credit — and only on the conditions you specify here.") { return "With a Creative Commons license, you keep your copyright but allow people to copy and distribute your work provided they give you credit — and only on the conditions you specify here."; } 
 if (s == "Taiwan") { return "Taiwan"; } 
 if (s == "If you desire a license governed by the Copyright Law of a specific jurisdiction, please select the appropriate jurisdiction.") { return "Om du önskar att din licens lyder under ett specifikt lands upphovsrättslagstiftning, var god välj lämplig jurisdiktion."; } 
 if (s == "Bulgaria") { return "Bulgarien"; } 
 if (s == "Romania") { return "Rumänien"; } 
 if (s == "Licensor permits others to make derivative works") { return "Licensor permits others to make derivative works"; } 
 if (s == "Portugal") { return "Portugal"; } 
 if (s == "Mexico") { return "Mexiko"; } 
 if (s == "work") { return "verk"; } 
 if (s == "India") { return "Indien"; } 
 if (s == "China Mainland") { return "Kina"; } 
 if (s == "Malaysia") { return "Malaysia"; } 
 if (s == "Austria") { return "Österrike"; } 
 if (s == "Colombia") { return "Columbia"; } 
 if (s == "Greece") { return "Grekland"; } 
 if (s == "Hungary") { return "Ungern"; } 
 if (s == "Share Alike") { return "Dela Lika"; } 
 if (s == "The licensor permits others to distribute derivative works only under the same license or one compatible with the one that governs the licensor's work.") { return "Licensgivaren tillåter andra att distribuera bearbetningar av verket endast under en licens som är identisk med den som gäller för licensgivarens verk."; } 
alert("Falling off the end.");
return s;
		}