var in_string = "<div id=\"cc_js_generated_box\">\n<div id=\"cc_js_lic-menu\">\n\n  <div id=\"cc_js_want_cc_license_at_all\">\n    <span>\n      <input checked=\"checked\" id=\"cc_js_want_cc_license_sure\" name=\"cc_js_want_cc_license\" onclick=\"cc_js_enable_widget();\" type=\"radio\" value=\"sure\"/><label class=\"cc_js_infobox\" for=\"cc_js_want_cc_license_sure\"><span onmouseout=\"cc_js_hide_tip()\" onmouseover=\"cc_js_on_tooltip_html(event,'&lt;p&gt;&lt;strong&gt;' + cc_js_t('Creative Commons') + '&lt;/strong&gt; ' + cc_js_t('With a Creative Commons license, you keep your copyright but allow people to copy and distribute your work provided they give you credit — and only on the conditions you specify here.') + '&lt;/p&gt;');\">A <span class=\"cc_js_question\">Creative Commons</span> license</span></label>\n    </span>\n    <span>\n\t    <input id=\"cc_js_want_cc_license_nah\" name=\"cc_js_want_cc_license\" onclick=\"cc_js_disable_widget();\" type=\"radio\" value=\"nah\"/>\n\t    <label for=\"cc_js_want_cc_license_nah\"><span>No license</span></label>\n    </span>\n  </div>\n\n  <div id=\"cc_js_required\">\n    \n    <p class=\"cc_js_hidden\">\n      <input checked=\"checked\" id=\"cc_js_share\" name=\"cc_js_share\" style=\"display: none;\" type=\"checkbox\" value=\"1\"/>\n    </p>\n      \n      \n    <p>\n      <input id=\"cc_js_remix\" name=\"cc_js_remix\" onclick=\"cc_js_modify(this);\" type=\"checkbox\" value=\"\"/>\n      <label class=\"cc_js_question\" for=\"cc_js_remix\" id=\"cc_js_remix-label\" onclick=\"cc_js_call_me_on_label_selection(this);\" onmouseout=\"cc_js_hide_tip()\" onmouseover=\"cc_js_on_tooltip_html(event,'&lt;p&gt;&lt;strong&gt;' + cc_js_t('Remix') + '&lt;/strong&gt; ' + cc_js_t('Licensor permits others to make derivative works') + '&lt;/p&gt;');\" style=\"color: black;\"><strong><span>Allow Remixing</span></strong></label> \n    </p>\n    \n    \n    <p>\n      <input id=\"cc_js_nc\" name=\"cc_js_nc\" onclick=\"cc_js_modify(this);\" type=\"checkbox\" value=\"\"/>\n      <label class=\"cc_js_question\" for=\"cc_js_nc\" id=\"cc_js_nc-label\" onclick=\"cc_js_call_me_on_label_selection(this);\" onmouseout=\"cc_js_hide_tip()\" onmouseover=\"cc_js_on_tooltip_html(event,'&lt;p&gt;&lt;img src=&quot;http://creativecommons.org/icon/nc/standard.gif&quot; alt=&quot;nc&quot; class=&quot;cc_js_icon&quot; /&gt;&lt;strong&gt;' + cc_js_t('Noncommercial') + '&lt;/strong&gt; ' + cc_js_t('The licensor permits others to copy, distribute and transmit the work. In return, licensees may not use the work for commercial purposes — unless they get the licensor\\'s permission.') + '&lt;/p&gt;');\" style=\"color: black;\"><strong><span>Prohibit Commercial Use</span></strong></label> \n    </p>\n\n    <p>\n      <input id=\"cc_js_sa\" name=\"cc_js_sa\" onclick=\"cc_js_modify(this);\" type=\"checkbox\" value=\"\"/>\n      <label class=\"cc_js_question\" for=\"cc_js_sa\" id=\"cc_js_sa-label\" onclick=\"cc_js_call_me_on_label_selection(this);\" onmouseout=\"cc_js_hide_tip()\" onmouseover=\"cc_js_on_tooltip_html(event,'&lt;p&gt;&lt;img src=&quot;http://creativecommons.org/icon/sa/standard.gif&quot; alt=&quot;sa&quot; class=&quot;cc_js_icon&quot; /&gt;&lt;strong&gt;' + cc_js_t('Share Alike') + '&lt;/strong&gt; ' + cc_js_t('The licensor permits others to distribute derivative works only under the same license or one compatible with the one that governs the licensor\\'s work.') + '&lt;/p&gt;');\" style=\"color: black;\"><strong><span>Require Share-Alike</span></strong></label>\n    </p>\n        \n    <br/>\n    \n    \n    \n  </div>\n  \n  <div id=\"cc_js_jurisdiction_box\">\n    <p><strong class=\"cc_js_question\" onmouseout=\"cc_js_hide_tip()\" onmouseover=\"cc_js_on_tooltip_html(event,'&lt;p&gt;&lt;strong&gt;Jurisdiction&lt;/strong&gt; ' + cc_js_t('If you desire a license governed by the Copyright Law of a specific jurisdiction, please select the appropriate jurisdiction.') + '&lt;/p&gt;');\"><span>Licensens jurisdiktion:</span></strong>  </p>\n    <select id=\"cc_js_jurisdiction\" name=\"cc_js_jurisdiction\" onchange=\"cc_js_modify(this);\" onclick=\"cc_js_modify(this);\">\n      \n      <option id=\"cc_js_jurisdiction_choice_generic\" value=\"generic\">Unported</option><option id=\"cc_js_jurisdiction_choice_ar\" value=\"ar\">Argentina</option><option id=\"cc_js_jurisdiction_choice_au\" value=\"au\">Australien</option><option id=\"cc_js_jurisdiction_choice_at\" value=\"at\">Österrike</option><option id=\"cc_js_jurisdiction_choice_be\" value=\"be\">Belgien</option><option id=\"cc_js_jurisdiction_choice_br\" value=\"br\">Brasilien</option><option id=\"cc_js_jurisdiction_choice_bg\" value=\"bg\">Bulgarien</option><option id=\"cc_js_jurisdiction_choice_ca\" value=\"ca\">Kanada</option><option id=\"cc_js_jurisdiction_choice_cl\" value=\"cl\">Chile</option><option id=\"cc_js_jurisdiction_choice_cn\" value=\"cn\">Kina</option><option id=\"cc_js_jurisdiction_choice_co\" value=\"co\">Columbia</option><option id=\"cc_js_jurisdiction_choice_hr\" value=\"hr\">Kroatien</option><option id=\"cc_js_jurisdiction_choice_hu\" value=\"hu\">Ungern</option><option id=\"cc_js_jurisdiction_choice_dk\" value=\"dk\">Danmark</option><option id=\"cc_js_jurisdiction_choice_fi\" value=\"fi\">Finland</option><option id=\"cc_js_jurisdiction_choice_fr\" value=\"fr\">Frankrike</option><option id=\"cc_js_jurisdiction_choice_de\" value=\"de\">Tyskland</option><option id=\"cc_js_jurisdiction_choice_il\" value=\"il\">Israel</option><option id=\"cc_js_jurisdiction_choice_in\" value=\"in\">Indien</option><option id=\"cc_js_jurisdiction_choice_it\" value=\"it\">Italien</option><option id=\"cc_js_jurisdiction_choice_jp\" value=\"jp\">Japan</option><option id=\"cc_js_jurisdiction_choice_kr\" value=\"kr\">Korea</option><option id=\"cc_js_jurisdiction_choice_mk\" value=\"mk\">Makedonien</option><option id=\"cc_js_jurisdiction_choice_my\" value=\"my\">Malaysia</option><option id=\"cc_js_jurisdiction_choice_mt\" value=\"mt\">Malta</option><option id=\"cc_js_jurisdiction_choice_mx\" value=\"mx\">Mexiko</option><option id=\"cc_js_jurisdiction_choice_nl\" value=\"nl\">Nederländerna</option><option id=\"cc_js_jurisdiction_choice_pe\" value=\"pe\">Peru</option><option id=\"cc_js_jurisdiction_choice_ph\" value=\"ph\">Filippinerna</option><option id=\"cc_js_jurisdiction_choice_pl\" value=\"pl\">Polen</option><option id=\"cc_js_jurisdiction_choice_pt\" value=\"pt\">Portugal</option><option id=\"cc_js_jurisdiction_choice_si\" value=\"si\">Slovenien</option><option id=\"cc_js_jurisdiction_choice_za\" value=\"za\">Sydafrika</option><option id=\"cc_js_jurisdiction_choice_es\" value=\"es\">Spanien</option><option id=\"cc_js_jurisdiction_choice_se\" value=\"se\">Sverige</option><option id=\"cc_js_jurisdiction_choice_ch\" value=\"ch\">Schweiz</option><option id=\"cc_js_jurisdiction_choice_tw\" value=\"tw\">Taiwan</option><option id=\"cc_js_jurisdiction_choice_uk\" value=\"uk\">UK: England &amp; Wales</option><option id=\"cc_js_jurisdiction_choice_scotland\" value=\"scotland\">UK: Skottland</option><option id=\"cc_js_jurisdiction_choice_us\" value=\"us\">Förenta Staterna</option><option id=\"cc_js_jurisdiction_choice_gr\" value=\"gr\">Grekland</option><option id=\"cc_js_jurisdiction_choice_lu\" value=\"lu\">Luxemburg</option><option id=\"cc_js_jurisdiction_choice_hk\" value=\"hk\">Hong Kong</option><option id=\"cc_js_jurisdiction_choice_nz\" value=\"nz\">Nya Zeeland</option><option id=\"cc_js_jurisdiction_choice_rs\" value=\"rs\">Serbien</option><option id=\"cc_js_jurisdiction_choice_pr\" value=\"pr\">Puerto Rico</option><option id=\"cc_js_jurisdiction_choice_ec\" value=\"ec\">Ecuador</option><option id=\"cc_js_jurisdiction_choice_no\" value=\"no\">Norway</option><option id=\"cc_js_jurisdiction_choice_sg\" value=\"sg\">Singapore</option><option id=\"cc_js_jurisdiction_choice_ro\" value=\"ro\">Rumänien</option><option id=\"cc_js_jurisdiction_choice_gt\" value=\"gt\">Guatemala</option><option id=\"cc_js_jurisdiction_choice_th\" value=\"th\">Thailand</option><option id=\"cc_js_jurisdiction_choice_cz\" value=\"cz\">Tjeckien</option>\n    </select>\n  </div>\n  \n  <div id=\"cc_js_license_selected\">\n    <div id=\"cc_js_license_example\"/>\n  </div>\n  \n  \n  <div id=\"cc_js_tip_cloak\" style=\"position:absolute; visibility:hidden; z-index:100\">hidden tip</div> \n</div>\n\n<form class=\"cc_js_hidden\" id=\"cc_js_cc_js_result_storage\">\n  <input id=\"cc_js_result_uri\" name=\"cc_js_result_uri\" type=\"hidden\" value=\"\"/>\n  <input id=\"cc_js_result_img\" name=\"cc_js_result_img\" type=\"hidden\" value=\"\"/>\n  <input id=\"cc_js_result_name\" name=\"cc_js_result_name\" type=\"hidden\" value=\"\"/>\n</form>\n  \n</div>";


var thisScript = /complete.js/;

var theScripts = document.getElementsByTagName('SCRIPT');

for (var i = 0 ; i < theScripts.length; i++) {

    if(theScripts[i].src.match(thisScript)) {

        var inForm = false;

        var currentNode = theScripts[i].parentNode;

        while (currentNode != null) {

            if (currentNode.nodeType == 1) {

                if (currentNode.tagName.toLowerCase() == 'form') {

                    inForm = true;

                    break;

                }

	    }

	    /* always */

	    currentNode = currentNode.parentNode;

        }

        

        if (inForm) {

	    /* if we are inside a form, we do not want to create

	       another form tag. So replace our FORM tag with

	       a DIV.

	    */

            in_string = in_string.replace('<form ', '<div ');

            in_string = in_string.replace('</form>', '</div>');

        }

        var my_div = document.createElement('DIV');

        my_div.innerHTML = in_string;



        theScripts[i].parentNode.insertBefore(my_div, theScripts[i]);

        theScripts[i].parentNode.removeChild(theScripts[i]);

	break;

    }

}
